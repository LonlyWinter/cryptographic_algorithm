`timescale 1ns/1ns

module test_uart;

reg clk;
reg rx;
reg tx;
reg status1;
reg status2;
reg status3;
reg status4;

serial_uart #(
    .CLK_FREQ(50),
    .BAUD(10)
) test_uart_inst (
    .clk(clk),
    .uart_rx(rx),
    .uart_tx(tx),
    .status1(status1),
    .status2(status2),
    .status3(status3),
    .status4(status4)
);

initial clk = 1;
always #2 clk = ~clk;

initial begin
    $dumpfile("test_uart.vcd");
    $dumpvars(0, test_uart);

    rx = 1;
    #52;

    // key = 64'h133457799BBCDFF1;
    // data_en = 64'h0123456789ABCDEF;
    // data_de = 64'h85E813540F0AB405;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    #2000;


    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    #2000;


    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    #2000;
    $finish;
end

endmodule
