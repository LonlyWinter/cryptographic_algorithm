`timescale 1ns/1ns

module test_uart;

reg clk;
reg rx;
reg tx;
reg status1;
reg status2;
reg status3;
reg status4;

serial_uart #(
    .CLK_FREQ(50),
    .BAUD(10)
) test_uart_inst (
    .clk(clk),
    .uart_rx(rx),
    .uart_tx(tx),
    .status1(status1),
    .status2(status2),
    .status3(status3),
    .status4(status4)
);

initial clk = 1;
always #2 clk = ~clk;

initial begin
    $dumpfile("test_uart.vcd");
    $dumpvars(0, test_uart);

    rx = 1;
    #52;

    // key = 64'h0123456789abcdef;
    // 00000001
    // 00100011
    // 010001010110011110001001101010111100110111101111
    // data_en = 64'h636f6d7075746572;
    // 0110001101101111011011010111000001110101011101000110010101110010
    // data_de = 64'h6a7d7274181d689f;
    // 0110101001111101011100100111010000011000000111010110100010011111
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    #100;


    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    #2000;


    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    rx = 1; #16;
    rx = 0; #16;
    rx = 1; #16;
    #2000;
    $finish;
end

endmodule
